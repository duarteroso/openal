module vopenal

//
pub struct AlcError {
pub mut:
	code int = 0
	msg  string = ''
}

pub fn alc_create_error(code int) AlcError {
	mut err := AlcError {
	}
	err.code = code
	err.msg = err.code_msg()
	return err
}

// code_str Return error code as string
pub fn (err &AlcError) code_str() string {
	return match err.code {
		alc_invalid_device		{ 'ALC_INVALID_DEVICE' }
		alc_invalid_context		{ 'ALC_INVALID_CONTEXT' }
		alc_invalid_enum 		{ 'ALC_INVALID_ENUM' }
		alc_invalid_value 		{ 'ALC_INVALID_VALUE' }
		alc_out_of_memory    	{ 'ALC_OUT_OF_MEMORY' }
		else					{ 'ALC_NO_ERROR' }
	}
}

// code_msg()
pub fn (err &AlcError) code_msg() string {
	return match err.code {
		alc_invalid_device		{ 'A bad device was passed to an OpenAL function' }
		alc_invalid_context 	{ 'A bad contet was passed to an OpenAL function' }
		alc_invalid_enum 		{ 'An unknown enum was passed to an OpenAL function' }
		alc_invalid_value 		{ 'An invalid value was passed to an OpenAL function' }
		alc_out_of_memory    	{ 'The requested operation resulted in OpenAL running out of memory' }
		else					{ 'There is not currently an error ' }
	}
}

// str Return error as string
pub fn (err &AlcError) str() string {
	return '${err.code_str()} - ${err.code_msg()}'
}