module vopenal

fn init() {
	//
}

// load_module loads OpenAL module
// Used to force the compiler to include the C pragmas
pub fn load_module() {
}

// unload_module unloads OpenAL module
pub fn unload_module() {
}
