module al

#flag linux -I/usr/include/AL
#flag linux -L/usr/lib64
#flag linux -lopenal

#include "AL/al.h"
