module al

type ALboolean = byte
type ALbooleanptr = voidptr

type ALchar = byte
type ALcharptr = charptr

type ALbyte = i8
type ALubyte = byte

type ALshort = i16
type ALushort = u16

type ALint = int
type ALintptr = voidptr

type ALuint = u32
type ALuintptr = voidptr

type ALsizei = int
type ALenum = int

type ALfloat = f32
type ALfloatptr = voidptr

type ALdouble = f64
type ALdoubleptr = voidptr
