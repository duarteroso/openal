module al

type ALboolean = byte
type ALchar = char
type ALbyte = i8
type ALubyte = byte
type ALshort = i16
type ALushort = u16
type ALint = int
type ALuint = u32
type ALsizei = int
type ALenum = int
type ALfloat = f32
type ALdouble = f64
