module al

type ALboolean = byte
type ALbooleanptr = &byte

type ALchar = byte
type ALcharptr = &char

type ALbyte = i8
type ALbyteptr = &i8

type ALubyte = byte
type ALubyteptr = &byte

type ALshort = i16
type ALushort = u16

type ALint = int
type ALintptr = &int

type ALuint = u32
type ALuintptr = &u32

type ALsizei = int
type ALenum = int

type ALfloat = f32
type ALfloatptr = &f32

type ALdouble = f64
type ALdoubleptr = &f64
