module al

fn C.alGetError() ALenum
