module alc

type ALCboolean = byte

type ALCchar = byte
type ALCcharptr = &char

type ALCbyte = i8
type ALCubyte = byte

type ALCshort = i16
type ALCushort = u16

type ALCint = int
type ALCintptr = &int

type ALCuint = u32

type ALCsizei = int

type ALCenum = int

type ALCfloat = f32

type ALCdouble = f64
