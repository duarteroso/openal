module al

// Runtime AL version
pub const (
	al_major_version = 1
	al_minor_version = 1
)

pub const (
	al_none  = 0
	al_false = 0
	al_true  = 1
)
