module alc

fn C.alcGetCurrentContext() &C.ALCcontext
