module al

fn C.alGetError() int
